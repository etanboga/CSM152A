`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:58:51 02/07/2019 
// Design Name: 
// Module Name:    Stopwatch_Top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Stopwatch_Top(
    );

Clock_Divider clk_div();
Seven_Seg_Controller disp(.digit0(), .digit1(), .digit2(), .digit3());

endmodule
